interface AdderInterface;
  logic [3:0] a, b;
  logic [4:0] sum;
endinterface
